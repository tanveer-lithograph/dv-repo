module testbench;
  initial begin
     $display("Hello asmicore");
     #1 $finish;
  end
endmodule
// let's start dv training
//no problem
// good commit
BUG_ON
// more changes
